`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 
// Design Name: 
// Module Name: W_Mem_2_4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`include "include.sv"

module W_Mem_2_4 #(parameter numWeight =30,
                             addressWidth = $clog2(numWeight), 
                             dataWidth = 16)
                             
                      ( 
                      input clk,
                      input wen,
                      input ren,
                      input [addressWidth-1:0] wadd,
                      input [addressWidth-1:0] radd,
                      input [dataWidth-1:0] win,
                      output logic [dataWidth-1:0] wout
                      );
        
    logic [dataWidth-1:0] mem [numWeight-1:0];
    
assign mem[0] =   16'b1111101010010001;
assign mem[1] =   16'b1111000011100111;
assign mem[2] =   16'b1111110111010000;
assign mem[3] =   16'b101001011010;
assign mem[4] =   16'b1101101110110;
assign mem[5] =   16'b1101111000100101;
assign mem[6] =   16'b111011111110;
assign mem[7] =   16'b1000010;
assign mem[8] =   16'b1111001011100111;
assign mem[9] =   16'b1110101011111000;
assign mem[10] =  16'b10110110101;
assign mem[11] =  16'b1111100011100001;
assign mem[12] =  16'b11000101111;
assign mem[13] =  16'b1111011111010101;
assign mem[14] =  16'b1111001101100101;
assign mem[15] =  16'b1010000100110;
assign mem[16] =  16'b110011101011;
assign mem[17] =  16'b101111011011;
assign mem[18] =  16'b110111000010;
assign mem[19] =  16'b1110101110110111;
assign mem[20] =  16'b1111101111001011;
assign mem[21] =  16'b1111011111110111;
assign mem[22] =  16'b1110101011110101;
assign mem[23] =  16'b1111101111101111;
assign mem[24] =  16'b100001111111;
assign mem[25] =  16'b1111001001011001;
assign mem[26] =  16'b101010100101;
assign mem[27] =  16'b10000110101;
assign mem[28] =  16'b1111001001010110;
assign mem[29] =  16'b101011001;
        

//		always_ff @(posedge clk)
//		begin
//			if (wen)
//			begin
//				mem[wadd] <= win;
//			end
			
//			else
//			begin
//			 //Do Nothing
//            end
//		end 

    
        always_ff @(posedge clk)
        begin
            if (ren)
            begin
                wout <= mem[radd];
            end
            
            else
            begin
             //Do Nothing
            end
        end 
endmodule