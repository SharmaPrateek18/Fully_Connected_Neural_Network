`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 
// Design Name: 
// Module Name: W_Mem_2_12
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`include "include.sv"

module W_Mem_2_12 #(parameter numWeight =30,
                             addressWidth = $clog2(numWeight), 
                             dataWidth = 16)
                             
                      ( 
                      input clk,
                      input wen,
                      input ren,
                      input [addressWidth-1:0] wadd,
                      input [addressWidth-1:0] radd,
                      input [dataWidth-1:0] win,
                      output logic [dataWidth-1:0] wout
                      );
        
    logic [dataWidth-1:0] mem [numWeight-1:0];
    
assign mem[0] =   16'b100011010110;
assign mem[1] =   16'b1010100010001;
assign mem[2] =   16'b11001010000;
assign mem[3] =   16'b1110110101111001;
assign mem[4] =   16'b1111110111111010;
assign mem[5] =   16'b1111011010011010;
assign mem[6] =   16'b101011010001;
assign mem[7] =   16'b1111100110101010;
assign mem[8] =   16'b11010000101;
assign mem[9] =   16'b1111100110;
assign mem[10] =  16'b1010010010010;
assign mem[11] =  16'b1111100000111011;
assign mem[12] =  16'b110010100;
assign mem[13] =  16'b1111100101100110;
assign mem[14] =  16'b1111101111111001;
assign mem[15] =  16'b100100001;
assign mem[16] =  16'b100010110110;
assign mem[17] =  16'b1110000000;
assign mem[18] =  16'b1111101011001000;
assign mem[19] =  16'b10111010001;
assign mem[20] =  16'b1111001000101101;
assign mem[21] =  16'b1110010110010001;
assign mem[22] =  16'b1111101111100101;
assign mem[23] =  16'b1000001000111;
assign mem[24] =  16'b1111111100111110;
assign mem[25] =  16'b110011000;
assign mem[26] =  16'b10110011110;
assign mem[27] =  16'b101101010110;
assign mem[28] =  16'b1111110100100110;
assign mem[29] =  16'b1111010000111001;
        

//		always_ff @(posedge clk)
//		begin
//			if (wen)
//			begin
//				mem[wadd] <= win;
//			end
			
//			else
//			begin
//			 //Do Nothing
//            end
//		end 

    
        always_ff @(posedge clk)
        begin
            if (ren)
            begin
                wout <= mem[radd];
            end
            
            else
            begin
             //Do Nothing
            end
        end 
endmodule