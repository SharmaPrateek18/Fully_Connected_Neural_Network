`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 
// Design Name: 
// Module Name: W_Mem_1_4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`include "include.sv"

module W_Mem_1_4 #(parameter numWeight =784,
                             addressWidth = $clog2(numWeight), 
                             dataWidth = 16)
                             
                      ( 
                      input clk,
                      input wen,
                      input ren,
                      input [addressWidth-1:0] wadd,
                      input [addressWidth-1:0] radd,
                      input [dataWidth-1:0] win,
                      output logic [dataWidth-1:0] wout
                      );
        
    logic [dataWidth-1:0] mem [numWeight-1:0];
    
assign mem[0] =   16'b1111111111110010;
assign mem[1] =   16'b101101;
assign mem[2] =   16'b1111111111101001;
assign mem[3] =   16'b1111111111010101;
assign mem[4] =   16'b1111111111000100;
assign mem[5] =   16'b10011;
assign mem[6] =   16'b1;
assign mem[7] =   16'b1111111111011111;
assign mem[8] =   16'b101;
assign mem[9] =   16'b101110;
assign mem[10] =  16'b1111111111010100;
assign mem[11] =  16'b1111111111010100;
assign mem[12] =  16'b1111111111100011;
assign mem[13] =  16'b1111111111010111;
assign mem[14] =  16'b111;
assign mem[15] =  16'b1011;
assign mem[16] =  16'b1111111111111000;
assign mem[17] =  16'b1111111111000110;
assign mem[18] =  16'b10100;
assign mem[19] =  16'b101;
assign mem[20] =  16'b10010;
assign mem[21] =  16'b0;
assign mem[22] =  16'b1111111111111111;
assign mem[23] =  16'b11111;
assign mem[24] =  16'b1111111111001110;
assign mem[25] =  16'b1010;
assign mem[26] =  16'b1101;
assign mem[27] =  16'b1011;
assign mem[28] =  16'b101000;
assign mem[29] =  16'b100;
assign mem[30] =  16'b1110;
assign mem[31] =  16'b1111111111101000;
assign mem[32] =  16'b11000;
assign mem[33] =  16'b11101;
assign mem[34] =  16'b1111111111111001;
assign mem[35] =  16'b110010;
assign mem[36] =  16'b111111;
assign mem[37] =  16'b10001;
assign mem[38] =  16'b1111111111101010;
assign mem[39] =  16'b1111111110111101;
assign mem[40] =  16'b10;
assign mem[41] =  16'b110011;
assign mem[42] =  16'b100;
assign mem[43] =  16'b1111111111110111;
assign mem[44] =  16'b1001010;
assign mem[45] =  16'b1111111111111100;
assign mem[46] =  16'b1111111111100110;
assign mem[47] =  16'b1111111111001101;
assign mem[48] =  16'b10010;
assign mem[49] =  16'b11001;
assign mem[50] =  16'b1111111111110100;
assign mem[51] =  16'b11110;
assign mem[52] =  16'b1000;
assign mem[53] =  16'b1010000;
assign mem[54] =  16'b111001;
assign mem[55] =  16'b110111;
assign mem[56] =  16'b11;
assign mem[57] =  16'b1111111111101111;
assign mem[58] =  16'b1010001;
assign mem[59] =  16'b11001;
assign mem[60] =  16'b1000110;
assign mem[61] =  16'b1111111111111011;
assign mem[62] =  16'b1111111110001110;
assign mem[63] =  16'b1111111110101001;
assign mem[64] =  16'b1111111110001001;
assign mem[65] =  16'b1111111100101110;
assign mem[66] =  16'b1111111011011000;
assign mem[67] =  16'b1111111010010100;
assign mem[68] =  16'b1111111010111010;
assign mem[69] =  16'b1111111010110100;
assign mem[70] =  16'b1111111011101000;
assign mem[71] =  16'b1111111011000000;
assign mem[72] =  16'b1111111100101100;
assign mem[73] =  16'b1111111011000101;
assign mem[74] =  16'b1111111101001010;
assign mem[75] =  16'b1111111011000001;
assign mem[76] =  16'b1111111011100111;
assign mem[77] =  16'b1111111011010101;
assign mem[78] =  16'b1111111101101101;
assign mem[79] =  16'b1111111110110110;
assign mem[80] =  16'b1101001;
assign mem[81] =  16'b1001001;
assign mem[82] =  16'b110;
assign mem[83] =  16'b1111111111011100;
assign mem[84] =  16'b1111111111110010;
assign mem[85] =  16'b11111;
assign mem[86] =  16'b1111111111100010;
assign mem[87] =  16'b1111111111110100;
assign mem[88] =  16'b1111111111010001;
assign mem[89] =  16'b1111111110110001;
assign mem[90] =  16'b1111111010111110;
assign mem[91] =  16'b1111111010111000;
assign mem[92] =  16'b1111111000011000;
assign mem[93] =  16'b1111111001011100;
assign mem[94] =  16'b1101000;
assign mem[95] =  16'b100110001;
assign mem[96] =  16'b1011;
assign mem[97] =  16'b1111111111100000;
assign mem[98] =  16'b1111111100110000;
assign mem[99] =  16'b1111111111001111;
assign mem[100] = 16'b1000001;
assign mem[101] = 16'b1011011000;
assign mem[102] = 16'b1001110101;
assign mem[103] = 16'b1111111111001011;
assign mem[104] = 16'b1111110100100000;
assign mem[105] = 16'b1111101110010101;
assign mem[106] = 16'b1111101110111011;
assign mem[107] = 16'b1111110011111101;
assign mem[108] = 16'b1111111010001001;
assign mem[109] = 16'b111001;
assign mem[110] = 16'b1111111111010110;
assign mem[111] = 16'b1111111111011011;
assign mem[112] = 16'b1111111111100101;
assign mem[113] = 16'b100010;
assign mem[114] = 16'b1111111111111101;
assign mem[115] = 16'b10100;
assign mem[116] = 16'b1111111110100110;
assign mem[117] = 16'b1111111111100011;
assign mem[118] = 16'b1111111011001111;
assign mem[119] = 16'b1111110101111111;
assign mem[120] = 16'b1111110101101011;
assign mem[121] = 16'b1111110101011111;
assign mem[122] = 16'b1111111100011110;
assign mem[123] = 16'b1000000101;
assign mem[124] = 16'b1111101110101011;
assign mem[125] = 16'b1111101001000011;
assign mem[126] = 16'b1111101001010010;
assign mem[127] = 16'b11010001;
assign mem[128] = 16'b111111000;
assign mem[129] = 16'b111000101;
assign mem[130] = 16'b100010011;
assign mem[131] = 16'b1111111100100001;
assign mem[132] = 16'b1111111101011101;
assign mem[133] = 16'b1111111011001010;
assign mem[134] = 16'b1111110011111010;
assign mem[135] = 16'b1111110110110101;
assign mem[136] = 16'b1111111111010100;
assign mem[137] = 16'b100000000;
assign mem[138] = 16'b10111000;
assign mem[139] = 16'b1111111111011100;
assign mem[140] = 16'b11100;
assign mem[141] = 16'b1111111111011001;
assign mem[142] = 16'b10011;
assign mem[143] = 16'b10001101;
assign mem[144] = 16'b1111111111010101;
assign mem[145] = 16'b1111110;
assign mem[146] = 16'b1111110111100101;
assign mem[147] = 16'b1111110100000001;
assign mem[148] = 16'b1111110110100000;
assign mem[149] = 16'b1111110100100111;
assign mem[150] = 16'b1111110010101100;
assign mem[151] = 16'b1111111111101000;
assign mem[152] = 16'b1111100101101000;
assign mem[153] = 16'b10111000100;
assign mem[154] = 16'b10101010000;
assign mem[155] = 16'b101111101011;
assign mem[156] = 16'b100100111001;
assign mem[157] = 16'b1100001001;
assign mem[158] = 16'b1111111101011001;
assign mem[159] = 16'b1111101110111001;
assign mem[160] = 16'b1111011110011000;
assign mem[161] = 16'b1111101101111001;
assign mem[162] = 16'b1111110111101001;
assign mem[163] = 16'b1111110101110011;
assign mem[164] = 16'b1111111001101111;
assign mem[165] = 16'b1101001;
assign mem[166] = 16'b1111111101111100;
assign mem[167] = 16'b1111111111000100;
assign mem[168] = 16'b1111111111110001;
assign mem[169] = 16'b1111111111110001;
assign mem[170] = 16'b110011;
assign mem[171] = 16'b1111111111100111;
assign mem[172] = 16'b111110;
assign mem[173] = 16'b111111110;
assign mem[174] = 16'b1111110111011000;
assign mem[175] = 16'b1111110001011010;
assign mem[176] = 16'b1111110111101001;
assign mem[177] = 16'b1111100110010011;
assign mem[178] = 16'b1000001011;
assign mem[179] = 16'b10001110;
assign mem[180] = 16'b1111110100100011;
assign mem[181] = 16'b11101010110;
assign mem[182] = 16'b100001110100;
assign mem[183] = 16'b1010001000001;
assign mem[184] = 16'b1001001000001;
assign mem[185] = 16'b100100100110;
assign mem[186] = 16'b1111110110001001;
assign mem[187] = 16'b1111101010001001;
assign mem[188] = 16'b1111110100100101;
assign mem[189] = 16'b1111110001000110;
assign mem[190] = 16'b1111111100110101;
assign mem[191] = 16'b1111110010010010;
assign mem[192] = 16'b1111110110110100;
assign mem[193] = 16'b1000111;
assign mem[194] = 16'b1111111100001100;
assign mem[195] = 16'b1111111101111100;
assign mem[196] = 16'b1111111111100101;
assign mem[197] = 16'b1001000;
assign mem[198] = 16'b110001;
assign mem[199] = 16'b11000101;
assign mem[200] = 16'b100011;
assign mem[201] = 16'b10;
assign mem[202] = 16'b1111110111111101;
assign mem[203] = 16'b1111110101110110;
assign mem[204] = 16'b1111101111010110;
assign mem[205] = 16'b1111110001100111;
assign mem[206] = 16'b1111110000011100;
assign mem[207] = 16'b1111100100010101;
assign mem[208] = 16'b1111011100000111;
assign mem[209] = 16'b1111111100111011;
assign mem[210] = 16'b101000010110;
assign mem[211] = 16'b1001110001000;
assign mem[212] = 16'b110000101111;
assign mem[213] = 16'b100101101;
assign mem[214] = 16'b1111111001110001;
assign mem[215] = 16'b1111100001111110;
assign mem[216] = 16'b1111111101110111;
assign mem[217] = 16'b1111111010101101;
assign mem[218] = 16'b1111110011110111;
assign mem[219] = 16'b1111111111001001;
assign mem[220] = 16'b1111111111001110;
assign mem[221] = 16'b101000110;
assign mem[222] = 16'b1111111101000000;
assign mem[223] = 16'b1111111111001000;
assign mem[224] = 16'b1111111111100110;
assign mem[225] = 16'b1110;
assign mem[226] = 16'b1010;
assign mem[227] = 16'b100011001;
assign mem[228] = 16'b100000111;
assign mem[229] = 16'b11011011;
assign mem[230] = 16'b1111111110101000;
assign mem[231] = 16'b1111111111111010;
assign mem[232] = 16'b1110011011;
assign mem[233] = 16'b1111111001111111;
assign mem[234] = 16'b1111111110100000;
assign mem[235] = 16'b1111110010001000;
assign mem[236] = 16'b1111101010111000;
assign mem[237] = 16'b1111111010011010;
assign mem[238] = 16'b1000010111110;
assign mem[239] = 16'b1010110110010;
assign mem[240] = 16'b10010001000;
assign mem[241] = 16'b1111110101011100;
assign mem[242] = 16'b1111111111011101;
assign mem[243] = 16'b101110;
assign mem[244] = 16'b1111111111011010;
assign mem[245] = 16'b1111111111111111;
assign mem[246] = 16'b1111111110101101;
assign mem[247] = 16'b10001101;
assign mem[248] = 16'b1111010011;
assign mem[249] = 16'b1000111110;
assign mem[250] = 16'b11111010;
assign mem[251] = 16'b100001;
assign mem[252] = 16'b100001;
assign mem[253] = 16'b101101;
assign mem[254] = 16'b1111111111111010;
assign mem[255] = 16'b101110001;
assign mem[256] = 16'b100111111;
assign mem[257] = 16'b1001000000;
assign mem[258] = 16'b101010011;
assign mem[259] = 16'b100011101010;
assign mem[260] = 16'b1001010011;
assign mem[261] = 16'b100100001;
assign mem[262] = 16'b11001011101;
assign mem[263] = 16'b1111110001001000;
assign mem[264] = 16'b1111011110100100;
assign mem[265] = 16'b1001111001;
assign mem[266] = 16'b1010001110011;
assign mem[267] = 16'b111110010001;
assign mem[268] = 16'b1111111100010010;
assign mem[269] = 16'b101000111;
assign mem[270] = 16'b110110010;
assign mem[271] = 16'b101101001;
assign mem[272] = 16'b1111111101001011;
assign mem[273] = 16'b1111111111010010;
assign mem[274] = 16'b1001110001;
assign mem[275] = 16'b10011010100;
assign mem[276] = 16'b1011001001;
assign mem[277] = 16'b1010111010;
assign mem[278] = 16'b111010011;
assign mem[279] = 16'b10000;
assign mem[280] = 16'b1111111110111011;
assign mem[281] = 16'b1111111111111111;
assign mem[282] = 16'b11110110;
assign mem[283] = 16'b111111100;
assign mem[284] = 16'b1010111010;
assign mem[285] = 16'b1111111001010111;
assign mem[286] = 16'b10110100010;
assign mem[287] = 16'b1011101101;
assign mem[288] = 16'b1111111011100000;
assign mem[289] = 16'b1111111111000010;
assign mem[290] = 16'b10011101011;
assign mem[291] = 16'b1111110011111111;
assign mem[292] = 16'b1111111001100010;
assign mem[293] = 16'b110100111000;
assign mem[294] = 16'b1011001100000;
assign mem[295] = 16'b100111011010;
assign mem[296] = 16'b1111111101101100;
assign mem[297] = 16'b10101110;
assign mem[298] = 16'b1111111101100111;
assign mem[299] = 16'b11100001;
assign mem[300] = 16'b1111111001100000;
assign mem[301] = 16'b11000001;
assign mem[302] = 16'b10001000101;
assign mem[303] = 16'b10110010101;
assign mem[304] = 16'b11100011;
assign mem[305] = 16'b1001101000;
assign mem[306] = 16'b110010110;
assign mem[307] = 16'b1111111110111010;
assign mem[308] = 16'b100111;
assign mem[309] = 16'b1111111111010111;
assign mem[310] = 16'b101010011;
assign mem[311] = 16'b101000110;
assign mem[312] = 16'b1110010000;
assign mem[313] = 16'b1111111100010101;
assign mem[314] = 16'b100010010111;
assign mem[315] = 16'b11010100000;
assign mem[316] = 16'b10001000110;
assign mem[317] = 16'b1100010110;
assign mem[318] = 16'b10110000110;
assign mem[319] = 16'b1010101001;
assign mem[320] = 16'b1111111001011001;
assign mem[321] = 16'b101000111001;
assign mem[322] = 16'b11100011001;
assign mem[323] = 16'b10100110101;
assign mem[324] = 16'b1111110100011111;
assign mem[325] = 16'b1010000101;
assign mem[326] = 16'b1111101101001111;
assign mem[327] = 16'b1111110111110000;
assign mem[328] = 16'b1111111100001101;
assign mem[329] = 16'b1111111011;
assign mem[330] = 16'b111001111;
assign mem[331] = 16'b1110011100;
assign mem[332] = 16'b1001010110;
assign mem[333] = 16'b1010110;
assign mem[334] = 16'b11111001;
assign mem[335] = 16'b1111111111111011;
assign mem[336] = 16'b1111111111110101;
assign mem[337] = 16'b11101;
assign mem[338] = 16'b1111101;
assign mem[339] = 16'b1100110;
assign mem[340] = 16'b10001011010;
assign mem[341] = 16'b100000111;
assign mem[342] = 16'b1001001011;
assign mem[343] = 16'b10000000001;
assign mem[344] = 16'b1111110110101110;
assign mem[345] = 16'b10010110110;
assign mem[346] = 16'b1111101111110010;
assign mem[347] = 16'b1111100010011111;
assign mem[348] = 16'b1111100111000101;
assign mem[349] = 16'b1111110110111110;
assign mem[350] = 16'b1111111010100001;
assign mem[351] = 16'b1111111101110011;
assign mem[352] = 16'b1111110101000100;
assign mem[353] = 16'b1000111001;
assign mem[354] = 16'b1111111111110001;
assign mem[355] = 16'b10000000010;
assign mem[356] = 16'b1111111001001010;
assign mem[357] = 16'b1011011001;
assign mem[358] = 16'b1010010001;
assign mem[359] = 16'b10100100;
assign mem[360] = 16'b1010011;
assign mem[361] = 16'b10010111;
assign mem[362] = 16'b101100110;
assign mem[363] = 16'b1101010;
assign mem[364] = 16'b1111111111111010;
assign mem[365] = 16'b101101;
assign mem[366] = 16'b1010100;
assign mem[367] = 16'b11000011;
assign mem[368] = 16'b1011000010;
assign mem[369] = 16'b1111110101010011;
assign mem[370] = 16'b1111111001011110;
assign mem[371] = 16'b100;
assign mem[372] = 16'b1111001100011110;
assign mem[373] = 16'b1111111001000110;
assign mem[374] = 16'b1111100110100010;
assign mem[375] = 16'b1111111110000111;
assign mem[376] = 16'b100010;
assign mem[377] = 16'b1111110100011101;
assign mem[378] = 16'b1001010110;
assign mem[379] = 16'b1111111000011111;
assign mem[380] = 16'b1111111001000011;
assign mem[381] = 16'b1111111011110100;
assign mem[382] = 16'b1111000100;
assign mem[383] = 16'b10010000011;
assign mem[384] = 16'b111110000;
assign mem[385] = 16'b10011110;
assign mem[386] = 16'b1111100;
assign mem[387] = 16'b1111101110110010;
assign mem[388] = 16'b1111111010010100;
assign mem[389] = 16'b100000010;
assign mem[390] = 16'b11011000;
assign mem[391] = 16'b1111111110111011;
assign mem[392] = 16'b1001111;
assign mem[393] = 16'b110110;
assign mem[394] = 16'b1000110;
assign mem[395] = 16'b11000000;
assign mem[396] = 16'b1111111010001001;
assign mem[397] = 16'b1111011011011111;
assign mem[398] = 16'b1111110011000011;
assign mem[399] = 16'b1111111111010000;
assign mem[400] = 16'b1111111100110011;
assign mem[401] = 16'b1111110001101111;
assign mem[402] = 16'b1111111001111001;
assign mem[403] = 16'b1111110011100100;
assign mem[404] = 16'b1111111111011000;
assign mem[405] = 16'b1001001000;
assign mem[406] = 16'b1111110110101011;
assign mem[407] = 16'b1111110100000000;
assign mem[408] = 16'b1111110111011100;
assign mem[409] = 16'b1111110000110001;
assign mem[410] = 16'b1111111011111010;
assign mem[411] = 16'b1111110011101010;
assign mem[412] = 16'b1111110101000010;
assign mem[413] = 16'b1111111110101011;
assign mem[414] = 16'b1111101111101101;
assign mem[415] = 16'b1111101010011101;
assign mem[416] = 16'b1111110111110110;
assign mem[417] = 16'b1111111110101000;
assign mem[418] = 16'b110001;
assign mem[419] = 16'b1111111111101011;
assign mem[420] = 16'b1111111111101010;
assign mem[421] = 16'b10100;
assign mem[422] = 16'b1001011;
assign mem[423] = 16'b1111111010111111;
assign mem[424] = 16'b1111111110110011;
assign mem[425] = 16'b10100010;
assign mem[426] = 16'b1111101100110100;
assign mem[427] = 16'b1111101000111001;
assign mem[428] = 16'b1111111101111010;
assign mem[429] = 16'b1111111100001000;
assign mem[430] = 16'b1111110000110100;
assign mem[431] = 16'b1111111100010101;
assign mem[432] = 16'b111101100;
assign mem[433] = 16'b100011010;
assign mem[434] = 16'b1111101110001010;
assign mem[435] = 16'b1111111110001011;
assign mem[436] = 16'b1111110100110011;
assign mem[437] = 16'b1111101111101110;
assign mem[438] = 16'b1111101011101000;
assign mem[439] = 16'b1111101101001110;
assign mem[440] = 16'b1111111101110101;
assign mem[441] = 16'b1111111110000011;
assign mem[442] = 16'b1111110000000011;
assign mem[443] = 16'b1111110010000101;
assign mem[444] = 16'b1100101;
assign mem[445] = 16'b1111111001111100;
assign mem[446] = 16'b1101110;
assign mem[447] = 16'b101100;
assign mem[448] = 16'b1111111111101010;
assign mem[449] = 16'b1010001;
assign mem[450] = 16'b101010;
assign mem[451] = 16'b1111111001011101;
assign mem[452] = 16'b100110001;
assign mem[453] = 16'b10010110111;
assign mem[454] = 16'b1111111100011010;
assign mem[455] = 16'b1111101110010111;
assign mem[456] = 16'b1111101110110111;
assign mem[457] = 16'b1111101010110110;
assign mem[458] = 16'b11001;
assign mem[459] = 16'b1111101011110111;
assign mem[460] = 16'b1111111011100010;
assign mem[461] = 16'b1001100110;
assign mem[462] = 16'b1111110001001001;
assign mem[463] = 16'b1111110000000101;
assign mem[464] = 16'b100010100;
assign mem[465] = 16'b10110111111;
assign mem[466] = 16'b1111111100000001;
assign mem[467] = 16'b1111110010000011;
assign mem[468] = 16'b1111110100100000;
assign mem[469] = 16'b1111011111001001;
assign mem[470] = 16'b1111111000010110;
assign mem[471] = 16'b1111110010001001;
assign mem[472] = 16'b1111111011110011;
assign mem[473] = 16'b1111111000100001;
assign mem[474] = 16'b1111111111111111;
assign mem[475] = 16'b1111111111110001;
assign mem[476] = 16'b1111111111100100;
assign mem[477] = 16'b1111111111101010;
assign mem[478] = 16'b1111111111001111;
assign mem[479] = 16'b1111111101001101;
assign mem[480] = 16'b10111100;
assign mem[481] = 16'b1101100101;
assign mem[482] = 16'b1111111001010110;
assign mem[483] = 16'b1111111101011001;
assign mem[484] = 16'b1101111;
assign mem[485] = 16'b1111110100010111;
assign mem[486] = 16'b1111111010011100;
assign mem[487] = 16'b1111110010000010;
assign mem[488] = 16'b110100101;
assign mem[489] = 16'b1100100011;
assign mem[490] = 16'b110111011;
assign mem[491] = 16'b1010110001;
assign mem[492] = 16'b10101011;
assign mem[493] = 16'b110010110;
assign mem[494] = 16'b1111111111010010;
assign mem[495] = 16'b1011101111;
assign mem[496] = 16'b1111110011000010;
assign mem[497] = 16'b1111011100101001;
assign mem[498] = 16'b1111101000111010;
assign mem[499] = 16'b1111110111100101;
assign mem[500] = 16'b1111111101010001;
assign mem[501] = 16'b1111111011101001;
assign mem[502] = 16'b1101;
assign mem[503] = 16'b1110111;
assign mem[504] = 16'b110001;
assign mem[505] = 16'b1;
assign mem[506] = 16'b1000001;
assign mem[507] = 16'b1111111001011100;
assign mem[508] = 16'b1111110111100000;
assign mem[509] = 16'b110010011;
assign mem[510] = 16'b1010010010;
assign mem[511] = 16'b1111101011011110;
assign mem[512] = 16'b1111100100011100;
assign mem[513] = 16'b1111110101101100;
assign mem[514] = 16'b111011110;
assign mem[515] = 16'b10010100101;
assign mem[516] = 16'b1111111110111101;
assign mem[517] = 16'b1111111100001111;
assign mem[518] = 16'b1111011111010001;
assign mem[519] = 16'b10001010001;
assign mem[520] = 16'b1110101;
assign mem[521] = 16'b1111110010100110;
assign mem[522] = 16'b1111111111101010;
assign mem[523] = 16'b111011101;
assign mem[524] = 16'b1111111110100001;
assign mem[525] = 16'b1111111011001011;
assign mem[526] = 16'b1111110111010101;
assign mem[527] = 16'b1111111010100010;
assign mem[528] = 16'b1111111001010001;
assign mem[529] = 16'b1111111100000111;
assign mem[530] = 16'b1000000;
assign mem[531] = 16'b111111;
assign mem[532] = 16'b1000011;
assign mem[533] = 16'b11;
assign mem[534] = 16'b11011111;
assign mem[535] = 16'b1111111100001000;
assign mem[536] = 16'b1111111110110101;
assign mem[537] = 16'b111000110;
assign mem[538] = 16'b1011001110;
assign mem[539] = 16'b1111101111011110;
assign mem[540] = 16'b1111101011111010;
assign mem[541] = 16'b1111101101111111;
assign mem[542] = 16'b110110010;
assign mem[543] = 16'b1111111111111100;
assign mem[544] = 16'b1011001111;
assign mem[545] = 16'b1111111101000011;
assign mem[546] = 16'b1111111111011100;
assign mem[547] = 16'b1111111111000011;
assign mem[548] = 16'b1110001101;
assign mem[549] = 16'b11101100;
assign mem[550] = 16'b1101110001;
assign mem[551] = 16'b1101010001;
assign mem[552] = 16'b1111111100100001;
assign mem[553] = 16'b1100011101;
assign mem[554] = 16'b111010101;
assign mem[555] = 16'b110010011;
assign mem[556] = 16'b10001010;
assign mem[557] = 16'b1110101;
assign mem[558] = 16'b111111;
assign mem[559] = 16'b10111;
assign mem[560] = 16'b10010;
assign mem[561] = 16'b1111111111011100;
assign mem[562] = 16'b101101;
assign mem[563] = 16'b1111111101110011;
assign mem[564] = 16'b1111111110011101;
assign mem[565] = 16'b1010010001;
assign mem[566] = 16'b10000110101;
assign mem[567] = 16'b1111110110000010;
assign mem[568] = 16'b1111110110110110;
assign mem[569] = 16'b1100101;
assign mem[570] = 16'b11000010;
assign mem[571] = 16'b10001111000;
assign mem[572] = 16'b1111111110100000;
assign mem[573] = 16'b0;
assign mem[574] = 16'b1010110011;
assign mem[575] = 16'b1111111110110001;
assign mem[576] = 16'b1111111001011111;
assign mem[577] = 16'b100011101;
assign mem[578] = 16'b1010000101;
assign mem[579] = 16'b10010010111;
assign mem[580] = 16'b101110011;
assign mem[581] = 16'b1000110111;
assign mem[582] = 16'b10000100110;
assign mem[583] = 16'b10000100100;
assign mem[584] = 16'b1000111011;
assign mem[585] = 16'b1000001000;
assign mem[586] = 16'b1011;
assign mem[587] = 16'b1111111111111001;
assign mem[588] = 16'b1111111111010000;
assign mem[589] = 16'b10;
assign mem[590] = 16'b111000;
assign mem[591] = 16'b1111111111000011;
assign mem[592] = 16'b1111111110110100;
assign mem[593] = 16'b1001001011;
assign mem[594] = 16'b1000100101;
assign mem[595] = 16'b1111111001101100;
assign mem[596] = 16'b1111101010000010;
assign mem[597] = 16'b1111111100110000;
assign mem[598] = 16'b111110001;
assign mem[599] = 16'b100100001;
assign mem[600] = 16'b11010;
assign mem[601] = 16'b1111110011011010;
assign mem[602] = 16'b1111111000100101;
assign mem[603] = 16'b1111111100110100;
assign mem[604] = 16'b1111111110011000;
assign mem[605] = 16'b1111111101000101;
assign mem[606] = 16'b110111111;
assign mem[607] = 16'b111111101;
assign mem[608] = 16'b1111111100110001;
assign mem[609] = 16'b1011110010;
assign mem[610] = 16'b1101110111;
assign mem[611] = 16'b100001110;
assign mem[612] = 16'b1100001111;
assign mem[613] = 16'b101011100;
assign mem[614] = 16'b1010;
assign mem[615] = 16'b11011;
assign mem[616] = 16'b10110;
assign mem[617] = 16'b0;
assign mem[618] = 16'b100111;
assign mem[619] = 16'b1111111111001100;
assign mem[620] = 16'b1111111110010111;
assign mem[621] = 16'b1111111111100001;
assign mem[622] = 16'b11110000;
assign mem[623] = 16'b100000100;
assign mem[624] = 16'b101111011;
assign mem[625] = 16'b1111111000100100;
assign mem[626] = 16'b1111110010011011;
assign mem[627] = 16'b1010110111;
assign mem[628] = 16'b1100000111;
assign mem[629] = 16'b1101010;
assign mem[630] = 16'b111100110;
assign mem[631] = 16'b1111111110011000;
assign mem[632] = 16'b111110111;
assign mem[633] = 16'b10010110000;
assign mem[634] = 16'b1100011011;
assign mem[635] = 16'b1111110011101000;
assign mem[636] = 16'b1111111011111011;
assign mem[637] = 16'b1001000010;
assign mem[638] = 16'b1100011011;
assign mem[639] = 16'b1010100110;
assign mem[640] = 16'b110011110;
assign mem[641] = 16'b11000;
assign mem[642] = 16'b1111111111100101;
assign mem[643] = 16'b10100;
assign mem[644] = 16'b1001010;
assign mem[645] = 16'b10010;
assign mem[646] = 16'b1111111111110111;
assign mem[647] = 16'b111110;
assign mem[648] = 16'b1111111110110110;
assign mem[649] = 16'b1111111110101011;
assign mem[650] = 16'b100110000;
assign mem[651] = 16'b110100111;
assign mem[652] = 16'b1111000001;
assign mem[653] = 16'b1101000011;
assign mem[654] = 16'b1011100;
assign mem[655] = 16'b10100011100;
assign mem[656] = 16'b10000010101;
assign mem[657] = 16'b11110010010;
assign mem[658] = 16'b1111100110;
assign mem[659] = 16'b10000101110;
assign mem[660] = 16'b111111010;
assign mem[661] = 16'b1111110001;
assign mem[662] = 16'b1111111100000111;
assign mem[663] = 16'b110000110;
assign mem[664] = 16'b10010100011;
assign mem[665] = 16'b1011100010;
assign mem[666] = 16'b1100111011;
assign mem[667] = 16'b1011011000;
assign mem[668] = 16'b1001101110;
assign mem[669] = 16'b1111111111111010;
assign mem[670] = 16'b1111111111011001;
assign mem[671] = 16'b11111;
assign mem[672] = 16'b1111111111110000;
assign mem[673] = 16'b1100;
assign mem[674] = 16'b1000110;
assign mem[675] = 16'b1010;
assign mem[676] = 16'b10001011;
assign mem[677] = 16'b1111111111111101;
assign mem[678] = 16'b10011100;
assign mem[679] = 16'b1001010;
assign mem[680] = 16'b10001000;
assign mem[681] = 16'b1110011;
assign mem[682] = 16'b11100100;
assign mem[683] = 16'b1111110110000010;
assign mem[684] = 16'b1111110110011101;
assign mem[685] = 16'b1111110011101001;
assign mem[686] = 16'b1110111;
assign mem[687] = 16'b111001110;
assign mem[688] = 16'b1111111000011111;
assign mem[689] = 16'b11111010;
assign mem[690] = 16'b11011000;
assign mem[691] = 16'b1110011011;
assign mem[692] = 16'b11010111000;
assign mem[693] = 16'b1011100011;
assign mem[694] = 16'b110101001;
assign mem[695] = 16'b110010010;
assign mem[696] = 16'b100100010;
assign mem[697] = 16'b111;
assign mem[698] = 16'b1111111111000010;
assign mem[699] = 16'b1111111111100010;
assign mem[700] = 16'b100;
assign mem[701] = 16'b1111111111101001;
assign mem[702] = 16'b1111111111110101;
assign mem[703] = 16'b101010;
assign mem[704] = 16'b1011001;
assign mem[705] = 16'b1011111;
assign mem[706] = 16'b100101100;
assign mem[707] = 16'b1100101111;
assign mem[708] = 16'b101110011;
assign mem[709] = 16'b101001110;
assign mem[710] = 16'b1111111111010111;
assign mem[711] = 16'b1111111101110001;
assign mem[712] = 16'b1111111110010000;
assign mem[713] = 16'b11001111;
assign mem[714] = 16'b1011000100;
assign mem[715] = 16'b1111110111111100;
assign mem[716] = 16'b1111110110100000;
assign mem[717] = 16'b1011110111;
assign mem[718] = 16'b111111100;
assign mem[719] = 16'b11110000110;
assign mem[720] = 16'b10101110110;
assign mem[721] = 16'b100000011;
assign mem[722] = 16'b10011001;
assign mem[723] = 16'b1111111100001101;
assign mem[724] = 16'b1111111111100001;
assign mem[725] = 16'b1111111111111111;
assign mem[726] = 16'b110011;
assign mem[727] = 16'b10011;
assign mem[728] = 16'b11011;
assign mem[729] = 16'b100001;
assign mem[730] = 16'b10101;
assign mem[731] = 16'b1111111110111111;
assign mem[732] = 16'b101110;
assign mem[733] = 16'b11000010;
assign mem[734] = 16'b10010101;
assign mem[735] = 16'b10101000;
assign mem[736] = 16'b1111111111010101;
assign mem[737] = 16'b1010010;
assign mem[738] = 16'b1011000000;
assign mem[739] = 16'b1111100101;
assign mem[740] = 16'b1101110101;
assign mem[741] = 16'b10000101111;
assign mem[742] = 16'b11010001001;
assign mem[743] = 16'b10010111000;
assign mem[744] = 16'b10101100000;
assign mem[745] = 16'b100000100;
assign mem[746] = 16'b1100001100;
assign mem[747] = 16'b1011001101;
assign mem[748] = 16'b110011000;
assign mem[749] = 16'b11010;
assign mem[750] = 16'b110;
assign mem[751] = 16'b1111111111101111;
assign mem[752] = 16'b10;
assign mem[753] = 16'b10101;
assign mem[754] = 16'b1111111111001010;
assign mem[755] = 16'b1111111111110000;
assign mem[756] = 16'b1111111111101100;
assign mem[757] = 16'b10000;
assign mem[758] = 16'b1100;
assign mem[759] = 16'b1111111111010100;
assign mem[760] = 16'b11110;
assign mem[761] = 16'b1101;
assign mem[762] = 16'b1000111;
assign mem[763] = 16'b11110101;
assign mem[764] = 16'b11100010;
assign mem[765] = 16'b111110;
assign mem[766] = 16'b10011;
assign mem[767] = 16'b1111111;
assign mem[768] = 16'b1100000;
assign mem[769] = 16'b111100;
assign mem[770] = 16'b1101100;
assign mem[771] = 16'b1010001;
assign mem[772] = 16'b111011;
assign mem[773] = 16'b1111111111011100;
assign mem[774] = 16'b10101;
assign mem[775] = 16'b1111;
assign mem[776] = 16'b10101;
assign mem[777] = 16'b1001111;
assign mem[778] = 16'b0;
assign mem[779] = 16'b1100;
assign mem[780] = 16'b1111111111001010;
assign mem[781] = 16'b100000;
assign mem[782] = 16'b110;
assign mem[783] = 16'b1111111111100110;
        

//		always_ff @(posedge clk)
//		begin
//			if (wen)
//			begin
//				mem[wadd] <= win;
//			end
			
//			else
//			begin
//			 //Do Nothing
//            end
//		end 

    
        always_ff @(posedge clk)
        begin
            if (ren)
            begin
                wout <= mem[radd];
            end
            
            else
            begin
             //Do Nothing
            end
        end 
endmodule